/****************************************************************************
 * rv_driver.svh
 ****************************************************************************/

/**
 * Class: rv_driver
 * 
 * TODO: Add class documentation
 */
class rv_driver #(int WIDTH=32) extends uvm_component;

	function new(string name, uvm_component parent);
		super.new(name, parent);
	endfunction


endclass


