/****************************************************************************
 * rv_agent_pkg.sv
 ****************************************************************************/
`include "uvm_macros.svh"

  
/**
 * Package: rv_agent_pkg
 * 
 * TODO: Add package documentation
 */
package rv_agent_pkg;
	import uvm_pkg::*;
	import tblink_rpc::*;
	
	`include "rv_initiator_agent.svh"
	`include "rv_initiator_bfm_impl.svh"
	`include "rv_initiator_driver.svh"


endpackage


