/****************************************************************************
 * rv_agent.svh
 ****************************************************************************/

  
/**
 * Class: rv_agent
 * 
 * TODO: Add class documentation
 */
class rv_agent #(int WIDTH=32) extends uvm_component;
	`uvm_component_utils(rv_agent)

	function new(string name, uvm_component parent);
		super.new(name, parent);
	endfunction
	
	function void build_phase(uvm_phase phase);
	endfunction


endclass


