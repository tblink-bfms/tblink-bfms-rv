/****************************************************************************
 * smoke_uvm_pkg.sv
 ****************************************************************************/
`include "uvm_macros.svh"

  
/**
 * Package: smoke_uvm_pkg
 * 
 * TODO: Add package documentation
 */
package smoke_uvm_pkg;
	import uvm_pkg::*;
	import tblink_rpc::*;
	import rv_agent_pkg::*;
	
	`include "smoke_uvm_test.svh"


endpackage


